[buckets]
0
[nodes]
)#���l֮R�I���볦�<�#������������̰� [nodes\]
137
[nodes]
)#���u�L<(j�'��FJG�9J            �� )#��,)Se��bڨK
��I�?�            {s [nodes\]
138
[nodes]
)#�y/x�����Ge��2ϓ�C�JN            � )#���#E��#�C�`}�ٓ;9z�             [nodes\]
139
[nodes]
)#�Ac����|=����L�p'm��            �i )#����볦�<�>�$^�/>>            U/ [nodes\]
140
[nodes]
)#��l֮R�I���볦�<�_w�            � )#�֮R�I���볦�<��_���            � )#����2�I.�W�QcY#5caMB�            ie )#��<�>�$^�G޳�m��V            �' )#��@�a;o`��d�>�U[]�V            � )#����yb��I��ǎD7ԣ��V            �� [nodes\]
141
[nodes]
)#���G��4�Ј)W���m���            T� )#��2j�*�t׈���� �_AX�            �� )#�($>42��{�H��IV��'�             ] )#�S�"<�Ds�j�o.�Ƃ,�o�F            9 )#��i�,7D��@|qC����            �e )#�0[�'a�|�P�3�]9 %T�            �� )#����!e��bj����3m�B            f� )#��#ZLe@j0�R/�QW��מ            {. [nodes\]
142
[nodes]
)#��hȀ?U�3�-1g��ѢO�v            � )#֟-z�%}^U�=�+ؚ��:�p�            � )#�礒��P&a�����_H)7            �� )#�%�#Y���jWBa��P�z            �� )#�s�������ώXX�3g��'            � )#�3��D5���?P�����=QI?            (� )#�k�7��o~z�AT8GM���            � )#�֮R�I���볦�<��S^<�            �� [nodes\]
143
[nodes]
)#T֮R�I���볦�<��w�G            {e )#z/&��~�@�����՝�
            7� )#MĿ)c	�ZCzoo����7I�            � [nodes\]
144
[nodes]
)"�Pup{ǘ��A%E���q�Sf�            � )"S����_c���wz��A�[��	            % )"�_�@�Ԣ�����a
v�\�"�            � )"�W�>a��9��܄���Z��            b� [nodes\]
145
[nodes]
)!���n�S�8FR��IZ�ƽ            �� ) ���>�2���Րr�>��oSR�            `� [nodes\]
146
[nodes]
)'ڥ(�:�`V�$rX _;��            � [nodes\]
147
[nodes]
),Rp�F�Ӳ^o&�i��g 7C��o            �� [nodes\]
149
[nodes]
)��G�- �Z
:�	�^��            57 [nodes\]
150
[nodes]
)YGjly9�¼���2�ì6H�]dC6            o� [nodes\]
152
[nodes]
(i�>
���y�ݓ�{���I��            C� [nodes\]
154
[nodes]
/�֣�`� +�����װ	��2N�K0            mb /�W$^�G޳M�C���>On��            �p -\���b���Qh./�	�Wm�            f� [nodes\]
156
[nodes]
< rsH���p���A8i�H!Wb�X������������� 2�NisQ�J�)ͺ����F|�gC��
������������� 7i`��F\�w�lO��A��E�o�            � 5.���\wZK��I��ֲGzl�b            �_ [nodes\]
157
[nodes]
 .Y.�]��\�r�r��2`m��	            	( uCy/!f�Z:�]�OJ@�m�Ms�            @ [nodes\]
158
[nodes]
B�PD�R�I���볦�<��^�Y            �B C��;�젞�c��iUu�	�.��j            h� A�0FBr��Au�����D*OeW�            �J F�<���I�r�2�9/�jU��s            mE GNj4�v��%��&�t�7�=ޙ            �G F,����G8S��jN�yPŗ�            �� E��
�>��{��[�0�<n�_�            �� @ 
��'��oͫ�������^	�            � [nodes\]
159
[nodes]
�!��ݔ����q��}7�x�(            w ƙ����K�arŘ��D*"�Q��            � ��wMyb�~��;���[��4��            ~� ���,��{���}^3��r�            �� ��$�:jTE�CT�e��1�Ú�H            �� �����3U��c�-E&�k�Qs�            \_ �<3��Q�����F��,1Yr-0            �� �?*�i9����CwI�O�{��]N�I            I� [nodes\]
[buckets\]
